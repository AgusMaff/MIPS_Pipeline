`timescale 1ns / 1ps

module ID_EX (
    input  wire        clk,
    input  wire        clk_en,        // Habilitar señal de reloj
    input  wire        reset,
    input  wire [31:0] id_dato_1,
    input  wire [31:0] id_dato_2,   
    input  wire [4:0]  id_rs,
    input  wire [4:0]  id_rt,
    input  wire [4:0]  id_rd,
    input  wire signed [31:0] id_extended_beq_offset,
    input  wire [5:0]  id_function_code,
    input  wire        id_ex_reg_dst,
    input  wire        id_ex_alu_src,
    input  wire [3:0]  id_ex_alu_op,
    input  wire        id_m_mem_read,
    input  wire        id_m_mem_write,
    input  wire        id_wb_mem_to_reg,
    input  wire        id_wb_reg_write,
    input  wire        id_ex_isJal,
    input  wire        id_ex_jalSel, // Bit de control para jalr
    input  wire [31:0] id_ex_pc_plus_8, // PC + 8 para la etapa ID/EX
    input  wire [2:0]  id_bhw_type,
    input  wire        id_ex_halt,
    input  wire        id_stall, 

    output reg [31:0] ex_dato_1,
    output reg [31:0] ex_dato_2,
    output reg [4:0]  ex_rs,
    output reg [4:0]  ex_rt,
    output reg [4:0]  ex_rd,
    output reg [5:0]  ex_function_code,
    output reg signed [31:0] ex_extended_beq_offset,
    output reg        ex_reg_dst,
    output reg        ex_alu_src,
    output reg [3:0]  ex_alu_op,
    output reg        ex_m_mem_read,
    output reg        ex_m_mem_write,
    output reg        ex_wb_mem_to_reg,
    output reg        ex_wb_reg_write,
    output reg        ex_isJal,
    output reg        ex_jalSel, // Bit de control para jalr
    output reg [31:0] ex_pc_plus_8, // PC + 8 para la etapa ID/EX
    output reg [2:0]  ex_bhw_type,
    output reg        ex_halt
);
    

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            ex_dato_1 <= 32'b0;
            ex_dato_2 <= 32'b0;
            ex_rs <= 5'b0;
            ex_rt <= 5'b0;
            ex_rd <= 5'b0;
            ex_function_code <= 6'b0;
            ex_extended_beq_offset <= 32'b0;
            ex_reg_dst <= 1'b0;
            ex_alu_src <= 1'b0;
            ex_alu_op <= 4'b0;
            ex_m_mem_read <= 1'b0;
            ex_m_mem_write <= 1'b0;
            ex_wb_mem_to_reg <= 1'b0;
            ex_wb_reg_write <= 1'b0;
            ex_bhw_type <= 3'b0;
            ex_halt <= 1'b0;
            ex_isJal <= 1'b0;
            ex_jalSel <= 1'b0; // Resetea el bit de control para jalr
            ex_pc_plus_8 <= 32'b0; // Resetea el PC + 8
        end 
        else if (id_stall && clk_en) begin
            // Inserta NOP en EX
            ex_dato_1 <= 32'b0;
            ex_dato_2 <= 32'b0;
            ex_rs <= 5'b0;
            ex_rt <= 5'b0;
            ex_rd <= 5'b0;
            ex_function_code <= 6'b0;
            ex_extended_beq_offset <= 32'b0;
            ex_reg_dst <= 1'b0;
            ex_alu_src <= 1'b0;
            ex_alu_op <= 4'b0;
            ex_m_mem_read <= 1'b0;
            ex_m_mem_write <= 1'b0;
            ex_wb_mem_to_reg <= 1'b0;
            ex_wb_reg_write <= 1'b0;
            ex_bhw_type <= 3'b0;
            ex_halt <= 1'b0;
            ex_isJal <= 1'b0;
            ex_jalSel <= 1'b0;
            ex_pc_plus_8 <= 32'b0;
        end 
        else if (clk_en) begin
            ex_dato_1 <= id_dato_1;
            ex_dato_2 <= id_dato_2;   
            ex_rs <= id_rs;
            ex_rt <= id_rt;
            ex_rd <= id_rd;
            ex_function_code <= id_function_code;
            ex_extended_beq_offset <= id_extended_beq_offset;
            ex_reg_dst <= id_ex_reg_dst;
            ex_alu_src <= id_ex_alu_src;
            ex_alu_op <= id_ex_alu_op;
            ex_m_mem_read <= id_m_mem_read;
            ex_m_mem_write <= id_m_mem_write;
            ex_wb_mem_to_reg <= id_wb_mem_to_reg;
            ex_wb_reg_write <= id_wb_reg_write; 
            ex_bhw_type <= id_bhw_type;
            ex_halt <= id_ex_halt;
            ex_isJal <= id_ex_isJal;
            ex_jalSel <= id_ex_jalSel; // Asigna el bit de control para jalr
            ex_pc_plus_8 <= id_ex_pc_plus_8;
        end
    end
endmodule